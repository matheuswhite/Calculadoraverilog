module OverflowDetection(A, B, Sum, Overflow);
	input A, B, Sum;
	output Overflow;
	
	
endmodule
